component pow_pll1 is
    port(outglobal_o: out std_logic;
         latch_i: in std_logic;
         outcore_o: out std_logic;
         ref_clk_i: in std_logic;
         rst_n_i: in std_logic);
end component;

__: pow_pll1 port map(outglobal_o=> , latch_i=> , outcore_o=> , ref_clk_i=> ,
    rst_n_i=> );